module dataDuplicator(input1, out1, out2);
	input [15:0] input1;
	output [15:0] out1, out2;
	
	assign out1 = input1;
	assign out2 = input1;
	
endmodule
